-Xshareclasses:none
